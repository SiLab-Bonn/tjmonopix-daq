//Verilog HDL for "TJ_Monopix_PADS", "decoupling_cap_filler" "functional"


module decoupling_cap_filler ( AVDD, AVSS, DVDD, DVSS, SUB );

  inout DVDD;
  inout AVSS;
  inout SUB;
  inout DVSS;
  inout AVDD;
endmodule

