//Verilog HDL for "pALPIDEfs_V2_BLOCKS_CAM", "PAD_PWELL" "functional"

`timescale 1ns / 1ps
module PAD_PWELL ( AVDD, AVSS, DVDD, DVSS, PWELL, SUB );

  inout PWELL;
  inout DVDD;
  inout AVSS;
  inout SUB;
  inout DVSS;
  inout AVDD;
endmodule
