//Verilog HDL for "TJ_Monopix_PADS", "PAD_ANALOG_IBIAS" "functional"


module PAD_ANALOG_IBIAS ( AVDD, AVSS, DVDD, DVSS, IBIAS, PAD, SUB );

  inout PAD;
  inout IBIAS;
  inout DVDD;
  inout AVSS;
  inout SUB;
  inout DVSS;
  inout AVDD;
endmodule
