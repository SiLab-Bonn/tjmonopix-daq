//Verilog HDL for "pALPIDEfs_V2_BLOCKS_CAM", "PAD_AVDD" "functional"
`timescale 1ns / 1ps

module PAD_AVDD ( AVDD, AVSS, DVDD, DVSS, SUB );

  inout DVDD;
  inout AVSS;
  inout SUB;
  inout DVSS;
  inout AVDD;
endmodule
