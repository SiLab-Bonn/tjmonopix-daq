//Verilog HDL for "pALPIDEfs_V2_BLOCKS_CAM", "PAD_SUB" "functional"


module PAD_SUB ( AVDD, AVSS, DVDD, DVSS, SUB );

  inout DVDD;
  inout AVSS;
  inout SUB;
  inout DVSS;
  inout AVDD;
endmodule
