//Verilog HDL for "TJ_Monopix_PADS", "PAD_ANALOG_NORES" "functional"


module PAD_ANALOG_NORES ( AVDD, AVSS, DVDD, DVSS, PAD, SUB );

  inout PAD;
  inout DVDD;
  inout AVSS;
  inout SUB;
  inout DVSS;
  inout AVDD;
endmodule
